library ieee;
use ieee.std_logic_1164.all;
 
entity de1_read is
    port(
        -- ADC
        ADC_CS_n : out std_logic;
        ADC_DIN  : out std_logic;
        ADC_DOUT : in  std_logic;
        ADC_SCLK : out std_logic;
      
        -- Audio
        AUD_ADCDAT  : in    std_logic;
        AUD_ADCLRCK : inout std_logic;
        AUD_BCLK    : inout std_logic;
        AUD_DACDAT  : out   std_logic;
        AUD_DACLRCK : inout std_logic;
        AUD_XCK     : out   std_logic;
      
        -- CLOCK
        CLOCK_50  : in std_logic;
        CLOCK2_50 : in std_logic;
        CLOCK3_50 : in std_logic;
        CLOCK4_50 : in std_logic;
      
        -- SDRAM
        DRAM_ADDR  : out   std_logic_vector(12 downto 0);
        DRAM_BA    : out   std_logic_vector(1 downto 0);
        DRAM_CAS_N : out   std_logic;
        DRAM_CKE   : out   std_logic;
        DRAM_CLK   : out   std_logic;
        DRAM_CS_N  : out   std_logic;
        DRAM_DQ    : inout std_logic_vector(15 downto 0);
        DRAM_LDQM  : out   std_logic;
        DRAM_RAS_N : out   std_logic;
        DRAM_UDQM  : out   std_logic;
        DRAM_WE_N  : out   std_logic;
      
        -- I2C for Audio and Video-In
        FPGA_I2C_SCLK : out   std_logic;
        FPGA_I2C_SDAT : inout std_logic;
      
        -- SEG7
        HEX0_N : out std_logic_vector(6 downto 0);
        HEX1_N : out std_logic_vector(6 downto 0);
        HEX2_N : out std_logic_vector(6 downto 0);
        HEX3_N : out std_logic_vector(6 downto 0);
        HEX4_N : out std_logic_vector(6 downto 0);
        HEX5_N : out std_logic_vector(6 downto 0);
      
        -- IR
        IRDA_RXD : in  std_logic;
        IRDA_TXD : out std_logic;
      
        -- KEY_N
        KEY_N : in std_logic_vector(3 downto 0);
      
        -- LED
        LEDR : out std_logic_vector(9 downto 0);
      
        -- PS2
        PS2_CLK  : inout std_logic;
        PS2_CLK2 : inout std_logic;
        PS2_DAT  : inout std_logic;
        PS2_DAT2 : inout std_logic;
      
        -- SW
        SW : in std_logic_vector(9 downto 0);
      
        -- Video-In
        TD_CLK27   : inout std_logic;
        TD_DATA    : out   std_logic_vector(7 downto 0);
        TD_HS      : out   std_logic;
        TD_RESET_N : out   std_logic;
        TD_VS      : out   std_logic;
      
        -- VGA
        VGA_B       : out std_logic_vector(7 downto 0);
        VGA_BLANK_N : out std_logic;
        VGA_CLK     : out std_logic;
        VGA_G       : out std_logic_vector(7 downto 0);
        VGA_HS      : out std_logic;
        VGA_R       : out std_logic_vector(7 downto 0);
        VGA_SYNC_N  : out std_logic;
        VGA_VS      : out std_logic;
      
        -- GPIO_0
        GPIO_0 : inout std_logic_vector(35 downto 0);
      
        -- GPIO_1
        GPIO_1 : inout std_logic_vector(35 downto 0)
          );         
end de1_read;
 
architecture rtl of de1_read is

	signal dbg_led_s 					: std_logic_vector(5 downto 0);
	signal stb_s						: std_logic_vector(5 downto 0);
	signal rxd_s						: std_logic_vector(5 downto 0);
	signal txd_s						: std_logic_vector(5 downto 0);
	
	signal frame_finished_s			: std_logic;
	signal sample_s					: std_logic;
	signal stuff_bit_s				: std_logic;
	signal bus_active_detect_s		: std_logic;
	signal rxd_sync_s					: std_logic;
	
	signal data_s						: std_logic_vector(63 downto 0);
	
	signal data_valid_s				: std_logic;

	signal uart_rxd : std_logic;
	signal uart_txd : std_logic;
begin

	stb_s <= "000000";


	shield_adapter_i0 : entity work.shield_adapter
		port map(
			gpio_b						=> GPIO_0,
			dbg_led_i					=> dbg_led_s,
			stb_i							=> stb_s,
			rxd_o							=> rxd_s,
			txd_i							=> txd_s
		);
		
	sampling_i0 : entity work.de1_sampling
		port map(
			clk							=> CLOCK_50,
			rst_n							=> KEY_N(0),
			
			rxd_i							=> rxd_s(0),
			frame_finished_i			=> frame_finished_s,
			
			rxd_sync_o					=> rxd_sync_s,
			sample_o						=> sample_s,
			stuff_bit_o					=> stuff_bit_s,
			bus_active_detect_o		=> bus_active_detect_s 
		);
		
	read_i0 : entity work.de1_core
		port map(
			clk							=> CLOCK_50,
			rst_n							=> KEY_N(0),
			
			rxd_sync_i					=> rxd_sync_s,
			sample_i						=> sample_s,
			stuff_bit_i					=> stuff_bit_s,
			bus_active_detect_i		=> bus_active_detect_s,
			
			frame_finished_o			=> frame_finished_s,
			
			data_o						=> data_s,
			valid_o						=> data_valid_s
		);
		
    debug_i0 : entity work.de1_debug
        generic map(
            widght_g                => 64
        )
        port map(
            clk                     => CLOCK_50,
            rst_n                   => KEY_N(0),

            data_i                  => data_s,
            valid_i                 => data_valid_s,

            rxd_i                   => uart_rxd,
            txd_o                   => uart_txd,
				GPIO_1						=> GPIO_1
        );
		  
		  GPIO_1(0) <= uart_rxd;
		  GPIO_1(1) <= uart_txd;
		  

		
	bin2hex_i0 : entity work.bin2hex
		port map(
			bin_i				=> data_s(3 downto 0),
			hex_o				=> HEX0_N
		);
		
	bin2hex_i1 : entity work.bin2hex
		port map(
			bin_i				=> data_s(7 downto 4),
			hex_o				=> HEX1_N
		);
		
	bin2hex_i2 : entity work.bin2hex
		port map(
			bin_i				=> data_s(11 downto 8),
			hex_o				=> HEX2_N
		);
		
	bin2hex_i3 : entity work.bin2hex
		port map(
			bin_i				=> data_s(15 downto 12),
			hex_o				=> HEX3_N
		);
		
	bin2hex_i4 : entity work.bin2hex
		port map(
			bin_i				=> data_s(19 downto 16),
			hex_o				=> HEX4_N
		);
		
	bin2hex_i5 : entity work.bin2hex
		port map(
			bin_i				=> data_s(23 downto 20),
			hex_o				=> HEX5_N
		);

end rtl;