library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity de1_sampling is
    port (
        clk                     : in    std_logic;
        rst_n                   : in    std_logic;

        rxd_i                   : in    std_logic;
        frame_finished_i        : in    std_logic;

        rxd_sync_o              : out   std_logic;
        sample_o                : out   std_logic;
        stuff_bit_o             : out   std_logic;
        bus_active_detect_o     : out   std_logic
    );
end entity;

architecture rtl of de1_sampling is

    signal rxd_async_s      : std_logic_vector(0 downto 0);
    signal rxd_sync_s       : std_logic_vector(0 downto 0);
    signal edge_s           : std_logic;
    signal sample_s         : std_logic;
    signal bus_active_s     : std_logic;
    signal stuff_bit_s      : std_logic;
    signal bit_stuff_error  : std_logic;
    signal hard_reload_s    : std_logic;
    signal sync_enable_s    : std_logic;

    signal rst_h            : std_logic;
begin
    rxd_async_s(0) <= rxd_i;
    rst_h  <= not rst_n;
    rxd_sync_o <= rxd_sync_s(0);
    sample_o <= sample_s;
    stuff_bit_o <= stuff_bit_s;
    bus_active_detect_o <= bus_active_s;

    sync_stage_i0 : entity work.olo_intf_sync
        generic map(
            RstLevel_g      => '1'
        )
        port map(
            Clk             => clk,
            Rst             => rst_h,
            DataAsync       => rxd_async_s,
            DataSync        => rxd_sync_s
        );

    edge_detect_i0 : entity work.edge_detect
        port map(
            clk             => clk,
            rst_n           => rst_n,

            data_i          => rxd_sync_s(0),

            edge_detect_o   => edge_s
        );

    sample_i0 : entity work.sample
        generic map(
            prescaler_g     => 4,
            sync_seg_g      => 1,
            prob_seg_g      => 5,
            phase_seg1_g    => 7,
            phase_seg2_g    => 7
        )
        port map(
            clk             => clk, 
            rst_n           => rst_n,

            edge_i        => edge_s,
            hard_reload_i   => hard_reload_s,
            sync_enable_i   => sync_enable_s,

            sample_o        => sample_s
        );

    idle_detect_i0 : entity work.idle_detect
        port map(
            clk             => clk,
            rst_n           => rst_n,

            frame_end_i     => frame_finished_i,
            edge_i          => edge_s,

            hard_reload_o   => hard_reload_s, 
            bus_active_o    => bus_active_s
        );

    destuffing_i0 : entity work.destuffing
        port map(
            clk             => clk,
            rst_n           => rst_n,

            data_i          => rxd_sync_s(0),
            sample_i        => sample_s,
            bus_active_i    => bus_active_s,
            
            stuff_bit_o     => stuff_bit_s,
            error_o          => bit_stuff_error
        );

    resync_validator_i0 : entity work.sample_validator
        port map(
            clk             => clk,
            rst_n           => rst_n,

            data_i          => rxd_sync_s(0),
            sample_i        => sample_s,
            edge_i          => edge_s,

            resync_valid_o  => sync_enable_s
        );



end architecture;